module Norgate(out, i1, i2);
    input i1, i2;
    output out;
    nor(out,i1,i2);
endmodule