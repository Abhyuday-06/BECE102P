module Andgate(out, i1, i2);
    input i1, i2;
    output out;
    and (out,i1,i2);
endmodule