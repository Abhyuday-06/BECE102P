module Xorgate(out, i1, i2);
    input i1, i2;
    output out;
    xor(out,i1,i2);
endmodule