module Nandgate(out, i1, i2);
    input i1, i2;
    output out;
    nand(out,i1,i2);
endmodule